module create_map(  
    input clk,
    input rst_sys,  
    input [1:0] state,
    input [4:0] num, //input num should be odd and between 3 and 19
    input [2:0] level,
    output reg [360:0] map
);  
integer i;
always @(posedge clk) begin
    if(state==2'b00)begin
    for(i = 0; i < 361; i = i + 1) begin
        map[i] = 1'b0;
    end
    if(level == 0&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 0&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=0;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=1;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 0&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=1;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 0&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=0;map[ 26]=0;map[ 27]=0;map[ 28]=0;map[ 29]=0;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=1;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=1;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=0;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=0;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=1;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=1;map[104]=1;map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 0&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=1;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=0;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=1;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=0;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;
        map[104]=0;map[105]=1;map[106]=0;map[107]=0;map[108]=0;map[109]=1;map[110]=0;map[111]=0;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=0;map[120]=1;map[121]=1;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;
        map[130]=0;map[131]=0;map[132]=0;map[133]=0;map[134]=0;map[135]=1;map[136]=0;map[137]=1;map[138]=0;map[139]=0;map[140]=0;map[141]=1;map[142]=0;
        map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=0;map[150]=1;map[151]=1;map[152]=1;map[153]=0;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 0&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=1;map[ 64]=0;map[ 65]=0;map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=0;map[ 96]=0;map[ 97]=0;map[ 98]=0;map[ 99]=0;map[100]=0;map[101]=1;map[102]=0;map[103]=0;map[104]=0;
        map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=1;map[114]=1;map[115]=1;map[116]=1;map[117]=1;map[118]=1;map[119]=0;
        map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=0;map[126]=0;map[127]=1;map[128]=0;map[129]=1;map[130]=0;map[131]=0;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=0;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=1;map[154]=0;map[155]=1;map[156]=0;map[157]=1;map[158]=0;map[159]=1;map[160]=0;map[161]=0;map[162]=0;map[163]=1;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=0;map[170]=1;map[171]=0;map[172]=1;map[173]=0;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=1;map[184]=0;map[185]=0;map[186]=0;map[187]=0;map[188]=0;map[189]=1;map[190]=0;map[191]=0;map[192]=0;map[193]=0;map[194]=0;
        map[195]=0;map[196]=1;map[197]=0;map[198]=1;map[199]=1;map[200]=1;map[201]=1;map[202]=1;map[203]=0;map[204]=1;map[205]=1;map[206]=1;map[207]=1;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 0&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=1;map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=1;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=1;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;
        map[102]=0;map[103]=0;map[104]=0;map[105]=0;map[106]=0;map[107]=1;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;
        map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;map[130]=1;map[131]=0;map[132]=1;map[133]=0;map[134]=1;map[135]=0;
        map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;map[143]=1;map[144]=0;map[145]=1;map[146]=0;map[147]=1;map[148]=0;map[149]=1;map[150]=0;map[151]=0;map[152]=0;
        map[153]=0;map[154]=1;map[155]=1;map[156]=1;map[157]=0;map[158]=1;map[159]=1;map[160]=1;map[161]=0;map[162]=1;map[163]=0;map[164]=1;map[165]=1;map[166]=1;map[167]=1;map[168]=1;map[169]=0;
        map[170]=0;map[171]=1;map[172]=0;map[173]=0;map[174]=0;map[175]=1;map[176]=0;map[177]=0;map[178]=0;map[179]=1;map[180]=0;map[181]=0;map[182]=0;map[183]=1;map[184]=0;map[185]=0;map[186]=0;
        map[187]=0;map[188]=1;map[189]=0;map[190]=1;map[191]=1;map[192]=1;map[193]=0;map[194]=1;map[195]=1;map[196]=1;map[197]=0;map[198]=1;map[199]=1;map[200]=1;map[201]=1;map[202]=1;map[203]=0;
        map[204]=0;map[205]=0;map[206]=0;map[207]=1;map[208]=0;map[209]=1;map[210]=0;map[211]=0;map[212]=0;map[213]=1;map[214]=0;map[215]=1;map[216]=0;map[217]=0;map[218]=0;map[219]=1;map[220]=0;
        map[221]=0;map[222]=1;map[223]=1;map[224]=1;map[225]=0;map[226]=1;map[227]=0;map[228]=1;map[229]=1;map[230]=1;map[231]=0;map[232]=1;map[233]=0;map[234]=1;map[235]=1;map[236]=1;map[237]=0;
        map[238]=0;map[239]=1;map[240]=0;map[241]=0;map[242]=0;map[243]=1;map[244]=0;map[245]=0;map[246]=0;map[247]=1;map[248]=0;map[249]=1;map[250]=0;map[251]=0;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=1;map[260]=1;map[261]=1;map[262]=1;map[263]=0;map[264]=1;map[265]=0;map[266]=1;map[267]=1;map[268]=1;map[269]=0;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 0&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=0;map[ 54]=0;map[ 55]=1;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=0;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=0;map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=1;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=1;map[110]=1;map[111]=0;map[112]=1;map[113]=0;
        map[114]=0;map[115]=0;map[116]=0;map[117]=1;map[118]=0;map[119]=1;map[120]=0;map[121]=0;map[122]=0;map[123]=0;map[124]=0;map[125]=1;map[126]=0;map[127]=1;map[128]=0;map[129]=0;map[130]=0;map[131]=1;map[132]=0;
        map[133]=0;map[134]=1;map[135]=1;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=0;map[142]=1;map[143]=1;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=0;map[150]=1;map[151]=0;
        map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=1;map[166]=0;map[167]=0;map[168]=0;map[169]=1;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=1;map[180]=1;map[181]=0;map[182]=1;map[183]=1;map[184]=1;map[185]=1;map[186]=1;map[187]=0;map[188]=1;map[189]=0;
        map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;map[195]=1;map[196]=0;map[197]=1;map[198]=0;map[199]=0;map[200]=0;map[201]=0;map[202]=0;map[203]=0;map[204]=0;map[205]=0;map[206]=0;map[207]=1;map[208]=0;
        map[209]=0;map[210]=1;map[211]=0;map[212]=1;map[213]=0;map[214]=1;map[215]=0;map[216]=1;map[217]=1;map[218]=1;map[219]=0;map[220]=1;map[221]=1;map[222]=1;map[223]=1;map[224]=1;map[225]=1;map[226]=1;map[227]=0;
        map[228]=0;map[229]=0;map[230]=0;map[231]=0;map[232]=0;map[233]=1;map[234]=0;map[235]=0;map[236]=0;map[237]=1;map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=0;map[244]=0;map[245]=1;map[246]=0;
        map[247]=0;map[248]=1;map[249]=1;map[250]=1;map[251]=1;map[252]=1;map[253]=0;map[254]=1;map[255]=1;map[256]=1;map[257]=1;map[258]=1;map[259]=0;map[260]=1;map[261]=0;map[262]=1;map[263]=0;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=1;map[270]=0;map[271]=1;map[272]=0;map[273]=1;map[274]=0;map[275]=1;map[276]=0;map[277]=1;map[278]=0;map[279]=0;map[280]=0;map[281]=1;map[282]=0;map[283]=1;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=0;map[290]=1;map[291]=0;map[292]=1;map[293]=0;map[294]=1;map[295]=0;map[296]=1;map[297]=0;map[298]=1;map[299]=1;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=1;map[306]=0;map[307]=1;map[308]=0;map[309]=0;map[310]=0;map[311]=1;map[312]=0;map[313]=0;map[314]=0;map[315]=1;map[316]=0;map[317]=0;map[318]=0;map[319]=1;map[320]=0;map[321]=1;map[322]=0;
        map[323]=0;map[324]=1;map[325]=0;map[326]=1;map[327]=0;map[328]=1;map[329]=1;map[330]=1;map[331]=0;map[332]=1;map[333]=1;map[334]=1;map[335]=1;map[336]=1;map[337]=0;map[338]=1;map[339]=0;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 1&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=1;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=0;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 1&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=0;map[ 18]=0;map[ 19]=1;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=0;map[ 32]=0;map[ 33]=1;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 1&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=1;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 1&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=0;map[ 26]=0;map[ 27]=0;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=1;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=0;map[ 52]=0;map[ 53]=0;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 1&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=0;map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=0;map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=1;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=1;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=0;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=1;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;
        map[104]=0;map[105]=1;map[106]=0;map[107]=1;map[108]=0;map[109]=0;map[110]=0;map[111]=1;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;
        map[130]=0;map[131]=1;map[132]=0;map[133]=1;map[134]=0;map[135]=1;map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;
        map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=0;map[150]=1;map[151]=0;map[152]=1;map[153]=1;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 1&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;map[ 65]=0;map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=1;map[ 98]=0;map[ 99]=0;map[100]=0;map[101]=0;map[102]=0;map[103]=1;map[104]=0;
        map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=0;map[112]=1;map[113]=1;map[114]=1;map[115]=0;map[116]=1;map[117]=1;map[118]=1;map[119]=0;
        map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=1;map[128]=0;map[129]=0;map[130]=0;map[131]=1;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=1;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=1;map[162]=0;map[163]=1;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=1;map[170]=1;map[171]=1;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=0;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=0;map[184]=0;map[185]=1;map[186]=0;map[187]=1;map[188]=0;map[189]=1;map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;
        map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=0;map[200]=1;map[201]=0;map[202]=1;map[203]=0;map[204]=1;map[205]=0;map[206]=1;map[207]=0;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 1&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=0;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=1;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=0;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=0;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=0;map[106]=0;map[107]=0;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;
        map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=1;map[124]=1;map[125]=1;map[126]=1;map[127]=0;map[128]=1;map[129]=1;map[130]=1;map[131]=1;map[132]=1;map[133]=0;map[134]=1;map[135]=0;
        map[136]=0;map[137]=0;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;map[143]=1;map[144]=0;map[145]=0;map[146]=0;map[147]=1;map[148]=0;map[149]=1;map[150]=0;map[151]=1;map[152]=0;
        map[153]=0;map[154]=1;map[155]=1;map[156]=1;map[157]=1;map[158]=1;map[159]=0;map[160]=1;map[161]=0;map[162]=1;map[163]=1;map[164]=1;map[165]=0;map[166]=1;map[167]=1;map[168]=1;map[169]=0;
        map[170]=0;map[171]=0;map[172]=0;map[173]=1;map[174]=0;map[175]=1;map[176]=0;map[177]=0;map[178]=0;map[179]=1;map[180]=0;map[181]=1;map[182]=0;map[183]=1;map[184]=0;map[185]=1;map[186]=0;
        map[187]=0;map[188]=1;map[189]=1;map[190]=1;map[191]=0;map[192]=1;map[193]=1;map[194]=1;map[195]=0;map[196]=1;map[197]=0;map[198]=1;map[199]=0;map[200]=1;map[201]=0;map[202]=1;map[203]=0;
        map[204]=0;map[205]=1;map[206]=0;map[207]=1;map[208]=0;map[209]=0;map[210]=0;map[211]=0;map[212]=0;map[213]=1;map[214]=0;map[215]=1;map[216]=0;map[217]=0;map[218]=0;map[219]=1;map[220]=0;
        map[221]=0;map[222]=1;map[223]=0;map[224]=1;map[225]=1;map[226]=1;map[227]=0;map[228]=1;map[229]=1;map[230]=1;map[231]=0;map[232]=1;map[233]=1;map[234]=1;map[235]=0;map[236]=1;map[237]=0;
        map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=0;map[246]=0;map[247]=1;map[248]=0;map[249]=0;map[250]=0;map[251]=1;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=0;map[257]=1;map[258]=1;map[259]=0;map[260]=1;map[261]=0;map[262]=1;map[263]=1;map[264]=1;map[265]=1;map[266]=1;map[267]=0;map[268]=1;map[269]=0;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 1&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=0;map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=1;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=0;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=0;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=0;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=1;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;
        map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;map[119]=1;map[120]=0;map[121]=0;map[122]=0;map[123]=1;map[124]=0;map[125]=0;map[126]=0;map[127]=0;map[128]=0;map[129]=0;map[130]=0;map[131]=1;map[132]=0;
        map[133]=0;map[134]=1;map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=1;map[150]=1;map[151]=0;
        map[152]=0;map[153]=0;map[154]=0;map[155]=1;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=1;map[162]=0;map[163]=1;map[164]=0;map[165]=1;map[166]=0;map[167]=1;map[168]=0;map[169]=1;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=1;map[176]=1;map[177]=1;map[178]=1;map[179]=0;map[180]=1;map[181]=0;map[182]=1;map[183]=0;map[184]=1;map[185]=0;map[186]=1;map[187]=0;map[188]=1;map[189]=0;
        map[190]=0;map[191]=0;map[192]=0;map[193]=0;map[194]=0;map[195]=1;map[196]=0;map[197]=1;map[198]=0;map[199]=0;map[200]=0;map[201]=1;map[202]=0;map[203]=0;map[204]=0;map[205]=1;map[206]=0;map[207]=1;map[208]=0;
        map[209]=0;map[210]=0;map[211]=0;map[212]=1;map[213]=1;map[214]=1;map[215]=0;map[216]=1;map[217]=0;map[218]=1;map[219]=1;map[220]=1;map[221]=1;map[222]=1;map[223]=0;map[224]=1;map[225]=0;map[226]=1;map[227]=0;
        map[228]=0;map[229]=1;map[230]=0;map[231]=0;map[232]=0;map[233]=1;map[234]=0;map[235]=1;map[236]=0;map[237]=1;map[238]=0;map[239]=1;map[240]=0;map[241]=0;map[242]=0;map[243]=1;map[244]=0;map[245]=1;map[246]=0;
        map[247]=0;map[248]=1;map[249]=1;map[250]=1;map[251]=1;map[252]=1;map[253]=0;map[254]=1;map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=1;map[260]=1;map[261]=0;map[262]=1;map[263]=0;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=1;map[270]=0;map[271]=1;map[272]=0;map[273]=0;map[274]=0;map[275]=1;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=1;map[282]=0;map[283]=0;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=0;map[290]=1;map[291]=1;map[292]=1;map[293]=0;map[294]=1;map[295]=1;map[296]=1;map[297]=1;map[298]=1;map[299]=0;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=0;map[306]=0;map[307]=0;map[308]=0;map[309]=1;map[310]=0;map[311]=1;map[312]=0;map[313]=0;map[314]=0;map[315]=0;map[316]=0;map[317]=1;map[318]=0;map[319]=0;map[320]=0;map[321]=1;map[322]=0;
        map[323]=0;map[324]=1;map[325]=1;map[326]=1;map[327]=1;map[328]=1;map[329]=0;map[330]=1;map[331]=1;map[332]=1;map[333]=1;map[334]=1;map[335]=0;map[336]=1;map[337]=0;map[338]=1;map[339]=1;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 2&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 2&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=1;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=0;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=0;map[ 39]=0;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 2&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=1;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 2&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=0;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 2&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=0;map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=1;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=1;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;
        map[104]=0;map[105]=0;map[106]=0;map[107]=1;map[108]=0;map[109]=0;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=1;map[120]=1;map[121]=1;map[122]=1;map[123]=0;map[124]=1;map[125]=0;map[126]=1;map[127]=1;map[128]=1;map[129]=0;
        map[130]=0;map[131]=1;map[132]=0;map[133]=0;map[134]=0;map[135]=0;map[136]=0;map[137]=1;map[138]=0;map[139]=0;map[140]=0;map[141]=1;map[142]=0;
        map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=0;map[150]=1;map[151]=1;map[152]=1;map[153]=0;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 2&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=1;map[ 64]=0;map[ 65]=0;map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=0;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;map[ 99]=1;map[100]=0;map[101]=1;map[102]=0;map[103]=1;map[104]=0;
        map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;map[114]=1;map[115]=0;map[116]=1;map[117]=0;map[118]=1;map[119]=0;
        map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=0;map[128]=0;map[129]=1;map[130]=0;map[131]=0;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=0;map[140]=1;map[141]=1;map[142]=1;map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=0;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=1;map[154]=0;map[155]=1;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=0;map[162]=0;map[163]=1;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=0;map[170]=1;map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=1;map[176]=1;map[177]=0;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=0;map[184]=0;map[185]=1;map[186]=0;map[187]=1;map[188]=0;map[189]=1;map[190]=0;map[191]=1;map[192]=0;map[193]=0;map[194]=0;
        map[195]=0;map[196]=1;map[197]=0;map[198]=1;map[199]=1;map[200]=1;map[201]=0;map[202]=1;map[203]=0;map[204]=1;map[205]=0;map[206]=1;map[207]=1;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 2&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=1;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=1;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=1;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=0;map[106]=0;map[107]=0;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=1;map[118]=0;
        map[119]=0;map[120]=1;map[121]=1;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;map[130]=1;map[131]=0;map[132]=1;map[133]=1;map[134]=1;map[135]=0;
        map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;map[143]=0;map[144]=0;map[145]=1;map[146]=0;map[147]=1;map[148]=0;map[149]=1;map[150]=0;map[151]=1;map[152]=0;
        map[153]=0;map[154]=1;map[155]=0;map[156]=1;map[157]=0;map[158]=1;map[159]=1;map[160]=1;map[161]=1;map[162]=1;map[163]=0;map[164]=1;map[165]=1;map[166]=1;map[167]=0;map[168]=1;map[169]=0;
        map[170]=0;map[171]=1;map[172]=0;map[173]=0;map[174]=0;map[175]=1;map[176]=0;map[177]=1;map[178]=0;map[179]=1;map[180]=0;map[181]=0;map[182]=0;map[183]=1;map[184]=0;map[185]=1;map[186]=0;
        map[187]=0;map[188]=1;map[189]=1;map[190]=1;map[191]=0;map[192]=1;map[193]=0;map[194]=1;map[195]=0;map[196]=1;map[197]=0;map[198]=1;map[199]=1;map[200]=1;map[201]=0;map[202]=1;map[203]=0;
        map[204]=0;map[205]=1;map[206]=0;map[207]=0;map[208]=0;map[209]=1;map[210]=0;map[211]=1;map[212]=0;map[213]=0;map[214]=0;map[215]=1;map[216]=0;map[217]=0;map[218]=0;map[219]=1;map[220]=0;
        map[221]=0;map[222]=1;map[223]=0;map[224]=1;map[225]=1;map[226]=1;map[227]=0;map[228]=1;map[229]=0;map[230]=1;map[231]=1;map[232]=1;map[233]=1;map[234]=1;map[235]=0;map[236]=1;map[237]=0;
        map[238]=0;map[239]=1;map[240]=0;map[241]=1;map[242]=0;map[243]=0;map[244]=0;map[245]=0;map[246]=0;map[247]=0;map[248]=0;map[249]=0;map[250]=0;map[251]=0;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=0;map[257]=0;map[258]=1;map[259]=1;map[260]=1;map[261]=1;map[262]=1;map[263]=1;map[264]=1;map[265]=1;map[266]=1;map[267]=0;map[268]=1;map[269]=1;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 2&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=0;map[ 50]=0;map[ 51]=0;map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=1;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=1;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=0;map[ 88]=0;map[ 89]=0;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=0;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=1;map[102]=1;map[103]=1;map[104]=1;map[105]=1;map[106]=1;map[107]=1;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;
        map[114]=0;map[115]=0;map[116]=0;map[117]=1;map[118]=0;map[119]=1;map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=1;map[128]=0;map[129]=1;map[130]=0;map[131]=0;map[132]=0;
        map[133]=0;map[134]=1;map[135]=1;map[136]=1;map[137]=0;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=1;map[148]=1;map[149]=1;map[150]=1;map[151]=0;
        map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=1;map[158]=0;map[159]=1;map[160]=0;map[161]=0;map[162]=0;map[163]=1;map[164]=0;map[165]=1;map[166]=0;map[167]=0;map[168]=0;map[169]=0;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=0;map[178]=1;map[179]=0;map[180]=1;map[181]=0;map[182]=1;map[183]=0;map[184]=1;map[185]=1;map[186]=1;map[187]=1;map[188]=1;map[189]=0;
        map[190]=0;map[191]=0;map[192]=0;map[193]=1;map[194]=0;map[195]=1;map[196]=0;map[197]=0;map[198]=0;map[199]=1;map[200]=0;map[201]=0;map[202]=0;map[203]=1;map[204]=0;map[205]=1;map[206]=0;map[207]=1;map[208]=0;
        map[209]=0;map[210]=1;map[211]=1;map[212]=1;map[213]=0;map[214]=1;map[215]=1;map[216]=1;map[217]=1;map[218]=1;map[219]=0;map[220]=1;map[221]=1;map[222]=1;map[223]=0;map[224]=1;map[225]=0;map[226]=1;map[227]=0;
        map[228]=0;map[229]=1;map[230]=0;map[231]=0;map[232]=0;map[233]=1;map[234]=0;map[235]=1;map[236]=0;map[237]=1;map[238]=0;map[239]=1;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=1;map[246]=0;
        map[247]=0;map[248]=1;map[249]=0;map[250]=1;map[251]=1;map[252]=1;map[253]=0;map[254]=1;map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=0;map[260]=1;map[261]=0;map[262]=1;map[263]=0;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=0;map[270]=0;map[271]=1;map[272]=0;map[273]=1;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=1;map[280]=0;map[281]=0;map[282]=0;map[283]=1;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=0;map[290]=0;map[291]=0;map[292]=1;map[293]=1;map[294]=1;map[295]=0;map[296]=1;map[297]=0;map[298]=1;map[299]=0;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=1;map[306]=0;map[307]=1;map[308]=0;map[309]=0;map[310]=0;map[311]=1;map[312]=0;map[313]=1;map[314]=0;map[315]=1;map[316]=0;map[317]=1;map[318]=0;map[319]=0;map[320]=0;map[321]=0;map[322]=0;
        map[323]=0;map[324]=1;map[325]=1;map[326]=1;map[327]=0;map[328]=1;map[329]=1;map[330]=1;map[331]=0;map[332]=1;map[333]=1;map[334]=1;map[335]=0;map[336]=1;map[337]=1;map[338]=1;map[339]=1;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 3&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 3&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=0;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;
        map[ 35]=0;map[ 36]=0;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 3&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=0;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=1;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 3&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=0;map[ 28]=0;map[ 29]=0;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=1;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=0;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=0;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=1;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=0;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 3&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=0;map[ 34]=0;map[ 35]=0;map[ 36]=0;map[ 37]=0;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=1;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=0;map[ 56]=0;map[ 57]=1;map[ 58]=0;map[ 59]=0;map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=1;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=1;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;
        map[104]=0;map[105]=1;map[106]=0;map[107]=1;map[108]=0;map[109]=0;map[110]=0;map[111]=0;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=0;map[120]=1;map[121]=1;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;
        map[130]=0;map[131]=0;map[132]=0;map[133]=1;map[134]=0;map[135]=1;map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;
        map[143]=0;map[144]=0;map[145]=1;map[146]=1;map[147]=0;map[148]=1;map[149]=0;map[150]=1;map[151]=0;map[152]=1;map[153]=1;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 3&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;map[ 65]=1;map[ 66]=0;map[ 67]=0;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=1;map[ 98]=0;map[ 99]=1;map[100]=0;map[101]=0;map[102]=0;map[103]=0;map[104]=0;
        map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;map[110]=1;map[111]=0;map[112]=1;map[113]=0;map[114]=1;map[115]=1;map[116]=1;map[117]=0;map[118]=1;map[119]=0;
        map[120]=0;map[121]=0;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=0;map[128]=0;map[129]=1;map[130]=0;map[131]=1;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=1;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=1;map[144]=1;map[145]=0;map[146]=1;map[147]=1;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=0;map[162]=0;map[163]=1;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=1;map[170]=1;map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=1;map[184]=0;map[185]=1;map[186]=0;map[187]=0;map[188]=0;map[189]=1;map[190]=0;map[191]=1;map[192]=0;map[193]=0;map[194]=0;
        map[195]=0;map[196]=0;map[197]=0;map[198]=1;map[199]=0;map[200]=1;map[201]=1;map[202]=1;map[203]=0;map[204]=1;map[205]=0;map[206]=1;map[207]=1;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 3&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=1;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=1;map[106]=0;map[107]=1;map[108]=0;map[109]=1;map[110]=0;map[111]=0;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;
        map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=0;map[124]=1;map[125]=0;map[126]=1;map[127]=1;map[128]=1;map[129]=0;map[130]=1;map[131]=0;map[132]=1;map[133]=0;map[134]=1;map[135]=0;
        map[136]=0;map[137]=1;map[138]=0;map[139]=0;map[140]=0;map[141]=0;map[142]=0;map[143]=1;map[144]=0;map[145]=0;map[146]=0;map[147]=1;map[148]=0;map[149]=1;map[150]=0;map[151]=1;map[152]=0;
        map[153]=0;map[154]=1;map[155]=1;map[156]=1;map[157]=0;map[158]=1;map[159]=1;map[160]=1;map[161]=0;map[162]=1;map[163]=1;map[164]=1;map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=0;
        map[170]=0;map[171]=1;map[172]=0;map[173]=1;map[174]=0;map[175]=1;map[176]=0;map[177]=1;map[178]=0;map[179]=0;map[180]=0;map[181]=1;map[182]=0;map[183]=1;map[184]=0;map[185]=0;map[186]=0;
        map[187]=0;map[188]=1;map[189]=0;map[190]=1;map[191]=0;map[192]=0;map[193]=0;map[194]=1;map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=0;map[200]=1;map[201]=1;map[202]=1;map[203]=0;
        map[204]=0;map[205]=0;map[206]=0;map[207]=1;map[208]=0;map[209]=0;map[210]=0;map[211]=1;map[212]=0;map[213]=0;map[214]=0;map[215]=1;map[216]=0;map[217]=1;map[218]=0;map[219]=1;map[220]=0;
        map[221]=0;map[222]=1;map[223]=1;map[224]=1;map[225]=0;map[226]=1;map[227]=0;map[228]=1;map[229]=1;map[230]=1;map[231]=0;map[232]=1;map[233]=0;map[234]=1;map[235]=0;map[236]=1;map[237]=0;
        map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=0;map[246]=0;map[247]=1;map[248]=0;map[249]=1;map[250]=0;map[251]=1;map[252]=0;map[253]=0;map[254]=0;
        map[255]=0;map[256]=1;map[257]=1;map[258]=1;map[259]=1;map[260]=1;map[261]=0;map[262]=0;map[263]=1;map[264]=1;map[265]=0;map[266]=1;map[267]=0;map[268]=1;map[269]=1;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 3&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=0;map[ 54]=0;map[ 55]=0;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=0;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=1;map[104]=1;map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;
        map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;map[119]=1;map[120]=0;map[121]=0;map[122]=0;map[123]=0;map[124]=0;map[125]=1;map[126]=0;map[127]=0;map[128]=0;map[129]=1;map[130]=0;map[131]=1;map[132]=0;
        map[133]=0;map[134]=1;map[135]=1;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=1;map[142]=1;map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=0;map[148]=1;map[149]=0;map[150]=1;map[151]=0;
        map[152]=0;map[153]=0;map[154]=0;map[155]=1;map[156]=0;map[157]=1;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=1;map[164]=0;map[165]=0;map[166]=0;map[167]=1;map[168]=0;map[169]=0;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;map[180]=1;map[181]=1;map[182]=1;map[183]=1;map[184]=1;map[185]=0;map[186]=1;map[187]=1;map[188]=1;map[189]=0;
        map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;map[195]=1;map[196]=0;map[197]=1;map[198]=0;map[199]=0;map[200]=0;map[201]=1;map[202]=0;map[203]=0;map[204]=0;map[205]=1;map[206]=0;map[207]=0;map[208]=0;
        map[209]=0;map[210]=1;map[211]=0;map[212]=1;map[213]=0;map[214]=1;map[215]=0;map[216]=1;map[217]=0;map[218]=1;map[219]=1;map[220]=1;map[221]=0;map[222]=1;map[223]=0;map[224]=1;map[225]=0;map[226]=1;map[227]=0;
        map[228]=0;map[229]=1;map[230]=0;map[231]=1;map[232]=0;map[233]=1;map[234]=0;map[235]=0;map[236]=0;map[237]=0;map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=0;map[244]=0;map[245]=1;map[246]=0;
        map[247]=0;map[248]=1;map[249]=0;map[250]=1;map[251]=0;map[252]=1;map[253]=1;map[254]=1;map[255]=1;map[256]=1;map[257]=1;map[258]=1;map[259]=1;map[260]=1;map[261]=1;map[262]=1;map[263]=1;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=1;map[270]=0;map[271]=0;map[272]=0;map[273]=1;map[274]=0;map[275]=1;map[276]=0;map[277]=1;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=1;map[290]=1;map[291]=0;map[292]=1;map[293]=0;map[294]=1;map[295]=0;map[296]=1;map[297]=1;map[298]=1;map[299]=1;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=1;map[306]=0;map[307]=1;map[308]=0;map[309]=0;map[310]=0;map[311]=1;map[312]=0;map[313]=0;map[314]=0;map[315]=1;map[316]=0;map[317]=1;map[318]=0;map[319]=1;map[320]=0;map[321]=0;map[322]=0;
        map[323]=0;map[324]=1;map[325]=0;map[326]=1;map[327]=0;map[328]=1;map[329]=1;map[330]=1;map[331]=0;map[332]=1;map[333]=1;map[334]=1;map[335]=0;map[336]=1;map[337]=0;map[338]=1;map[339]=1;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 4&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=1;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 4&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=0;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=0;map[ 32]=0;map[ 33]=0;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 4&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=1;map[ 66]=0;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 4&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=1;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=1;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=0;map[ 96]=0;map[ 97]=1;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 4&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=0;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=1;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=0;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;
        map[104]=0;map[105]=0;map[106]=0;map[107]=0;map[108]=0;map[109]=1;map[110]=0;map[111]=0;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=0;map[120]=1;map[121]=1;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;
        map[130]=0;map[131]=1;map[132]=0;map[133]=0;map[134]=0;map[135]=1;map[136]=0;map[137]=0;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;
        map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=1;map[150]=1;map[151]=0;map[152]=1;map[153]=1;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 4&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;map[ 65]=1;map[ 66]=0;map[ 67]=0;map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;map[ 99]=1;map[100]=0;map[101]=1;map[102]=0;map[103]=1;map[104]=0;
        map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;map[114]=1;map[115]=0;map[116]=1;map[117]=0;map[118]=1;map[119]=0;
        map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=0;map[128]=0;map[129]=1;map[130]=0;map[131]=0;map[132]=0;map[133]=0;map[134]=0;
        map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=1;map[144]=1;map[145]=1;map[146]=1;map[147]=1;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=0;map[154]=0;map[155]=0;map[156]=0;map[157]=1;map[158]=0;map[159]=0;map[160]=0;map[161]=1;map[162]=0;map[163]=0;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=1;map[170]=1;map[171]=1;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=0;map[184]=0;map[185]=0;map[186]=0;map[187]=0;map[188]=0;map[189]=1;map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;
        map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=0;map[200]=1;map[201]=1;map[202]=1;map[203]=1;map[204]=1;map[205]=0;map[206]=1;map[207]=0;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 4&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=1;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=1;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=1;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=0;map[106]=0;map[107]=0;map[108]=0;map[109]=0;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=1;map[116]=0;map[117]=0;map[118]=0;
        map[119]=0;map[120]=1;map[121]=1;map[122]=1;map[123]=1;map[124]=1;map[125]=1;map[126]=1;map[127]=0;map[128]=1;map[129]=1;map[130]=1;map[131]=0;map[132]=1;map[133]=0;map[134]=1;map[135]=0;
        map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;map[143]=1;map[144]=0;map[145]=0;map[146]=0;map[147]=1;map[148]=0;map[149]=0;map[150]=0;map[151]=1;map[152]=0;
        map[153]=0;map[154]=1;map[155]=0;map[156]=1;map[157]=0;map[158]=1;map[159]=1;map[160]=1;map[161]=0;map[162]=1;map[163]=1;map[164]=1;map[165]=1;map[166]=1;map[167]=1;map[168]=1;map[169]=0;
        map[170]=0;map[171]=1;map[172]=0;map[173]=0;map[174]=0;map[175]=0;map[176]=0;map[177]=1;map[178]=0;map[179]=0;map[180]=0;map[181]=0;map[182]=0;map[183]=1;map[184]=0;map[185]=0;map[186]=0;
        map[187]=0;map[188]=1;map[189]=1;map[190]=1;map[191]=1;map[192]=1;map[193]=0;map[194]=1;map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=1;map[200]=1;map[201]=1;map[202]=1;map[203]=0;
        map[204]=0;map[205]=1;map[206]=0;map[207]=1;map[208]=0;map[209]=1;map[210]=0;map[211]=1;map[212]=0;map[213]=0;map[214]=0;map[215]=1;map[216]=0;map[217]=1;map[218]=0;map[219]=0;map[220]=0;
        map[221]=0;map[222]=1;map[223]=0;map[224]=1;map[225]=0;map[226]=1;map[227]=0;map[228]=1;map[229]=1;map[230]=1;map[231]=0;map[232]=1;map[233]=0;map[234]=1;map[235]=0;map[236]=0;map[237]=0;
        map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=1;map[246]=0;map[247]=0;map[248]=0;map[249]=1;map[250]=0;map[251]=0;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=1;map[257]=1;map[258]=1;map[259]=0;map[260]=1;map[261]=0;map[262]=1;map[263]=0;map[264]=1;map[265]=1;map[266]=1;map[267]=1;map[268]=1;map[269]=1;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 4&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=1;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=0;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=0;map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=0;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=1;map[102]=1;map[103]=0;map[104]=1;map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;
        map[114]=0;map[115]=1;map[116]=0;map[117]=0;map[118]=0;map[119]=1;map[120]=0;map[121]=1;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=0;map[128]=0;map[129]=0;map[130]=0;map[131]=1;map[132]=0;
        map[133]=0;map[134]=1;map[135]=0;map[136]=1;map[137]=1;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=1;map[150]=1;map[151]=0;
        map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=1;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=1;map[166]=0;map[167]=0;map[168]=0;map[169]=1;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;map[180]=1;map[181]=1;map[182]=1;map[183]=1;map[184]=1;map[185]=1;map[186]=1;map[187]=1;map[188]=1;map[189]=0;
        map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;map[195]=0;map[196]=0;map[197]=1;map[198]=0;map[199]=0;map[200]=0;map[201]=1;map[202]=0;map[203]=0;map[204]=0;map[205]=1;map[206]=0;map[207]=0;map[208]=0;
        map[209]=0;map[210]=1;map[211]=0;map[212]=1;map[213]=1;map[214]=1;map[215]=0;map[216]=1;map[217]=0;map[218]=1;map[219]=1;map[220]=1;map[221]=1;map[222]=1;map[223]=0;map[224]=1;map[225]=1;map[226]=1;map[227]=0;
        map[228]=0;map[229]=1;map[230]=0;map[231]=1;map[232]=0;map[233]=1;map[234]=0;map[235]=1;map[236]=0;map[237]=1;map[238]=0;map[239]=1;map[240]=0;map[241]=0;map[242]=0;map[243]=0;map[244]=0;map[245]=1;map[246]=0;
        map[247]=0;map[248]=1;map[249]=0;map[250]=1;map[251]=0;map[252]=1;map[253]=0;map[254]=1;map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=1;map[260]=1;map[261]=0;map[262]=1;map[263]=1;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=0;map[270]=0;map[271]=0;map[272]=0;map[273]=1;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=1;map[282]=0;map[283]=1;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=0;map[290]=1;map[291]=1;map[292]=1;map[293]=1;map[294]=1;map[295]=1;map[296]=1;map[297]=0;map[298]=1;map[299]=1;map[300]=1;map[301]=0;map[302]=1;map[303]=0;
        map[304]=0;map[305]=1;map[306]=0;map[307]=1;map[308]=0;map[309]=1;map[310]=0;map[311]=1;map[312]=0;map[313]=0;map[314]=0;map[315]=1;map[316]=0;map[317]=1;map[318]=0;map[319]=1;map[320]=0;map[321]=0;map[322]=0;
        map[323]=0;map[324]=1;map[325]=1;map[326]=1;map[327]=0;map[328]=1;map[329]=0;map[330]=1;map[331]=1;map[332]=1;map[333]=0;map[334]=1;map[335]=0;map[336]=1;map[337]=0;map[338]=1;map[339]=1;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 5&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=1;map[ 14]=0;
        map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 5&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=0;map[ 18]=0;map[ 19]=0;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=0;map[ 32]=0;map[ 33]=0;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 5&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=0;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=0;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=0;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 5&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=0;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=0;map[ 52]=0;map[ 53]=1;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=1;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=0;map[ 96]=0;map[ 97]=1;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;map[104]=1;map[105]=1;map[106]=0;map[107]=0;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 5&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=0;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=0;map[ 56]=0;map[ 57]=1;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=0;map[ 62]=0;map[ 63]=1;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=0;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=1;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=1;map[102]=1;map[103]=0;
        map[104]=0;map[105]=1;map[106]=0;map[107]=1;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;
        map[117]=0;map[118]=1;map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=0;map[124]=1;map[125]=1;map[126]=1;map[127]=1;map[128]=1;map[129]=0;
        map[130]=0;map[131]=1;map[132]=0;map[133]=1;map[134]=0;map[135]=1;map[136]=0;map[137]=1;map[138]=0;map[139]=0;map[140]=0;map[141]=0;map[142]=0;
        map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=0;map[150]=1;map[151]=1;map[152]=1;map[153]=1;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 5&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;map[ 65]=0;map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=1;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;map[ 95]=0;map[ 96]=0;map[ 97]=1;map[ 98]=0;map[ 99]=0;map[100]=0;map[101]=1;map[102]=0;map[103]=1;map[104]=0;
        map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=0;map[114]=1;map[115]=1;map[116]=1;map[117]=0;map[118]=1;map[119]=0;
        map[120]=0;map[121]=0;map[122]=0;map[123]=1;map[124]=0;map[125]=1;map[126]=0;map[127]=1;map[128]=0;map[129]=1;map[130]=0;map[131]=0;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=1;map[138]=1;map[139]=0;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=1;map[146]=1;map[147]=0;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=1;map[154]=0;map[155]=0;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=1;map[162]=0;map[163]=0;map[164]=0;
        map[165]=0;map[166]=1;map[167]=0;map[168]=1;map[169]=0;map[170]=1;map[171]=1;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=0;map[178]=0;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=1;map[184]=0;map[185]=1;map[186]=0;map[187]=1;map[188]=0;map[189]=1;map[190]=0;map[191]=0;map[192]=0;map[193]=1;map[194]=0;
        map[195]=0;map[196]=1;map[197]=0;map[198]=1;map[199]=0;map[200]=1;map[201]=0;map[202]=1;map[203]=0;map[204]=1;map[205]=1;map[206]=1;map[207]=1;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 5&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=0;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=1;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=0;map[ 90]=1;map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=1;map[106]=0;map[107]=0;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;map[117]=0;map[118]=0;
        map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=1;map[124]=1;map[125]=0;map[126]=1;map[127]=0;map[128]=1;map[129]=0;map[130]=1;map[131]=0;map[132]=1;map[133]=0;map[134]=1;map[135]=0;
        map[136]=0;map[137]=0;map[138]=0;map[139]=1;map[140]=0;map[141]=1;map[142]=0;map[143]=1;map[144]=0;map[145]=1;map[146]=0;map[147]=0;map[148]=0;map[149]=0;map[150]=0;map[151]=1;map[152]=0;
        map[153]=0;map[154]=1;map[155]=1;map[156]=1;map[157]=0;map[158]=1;map[159]=0;map[160]=1;map[161]=0;map[162]=1;map[163]=1;map[164]=1;map[165]=1;map[166]=1;map[167]=1;map[168]=1;map[169]=0;
        map[170]=0;map[171]=1;map[172]=0;map[173]=1;map[174]=0;map[175]=1;map[176]=0;map[177]=1;map[178]=0;map[179]=0;map[180]=0;map[181]=1;map[182]=0;map[183]=0;map[184]=0;map[185]=1;map[186]=0;
        map[187]=0;map[188]=1;map[189]=0;map[190]=1;map[191]=0;map[192]=1;map[193]=0;map[194]=1;map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=1;map[200]=1;map[201]=0;map[202]=1;map[203]=0;
        map[204]=0;map[205]=0;map[206]=0;map[207]=1;map[208]=0;map[209]=1;map[210]=0;map[211]=1;map[212]=0;map[213]=0;map[214]=0;map[215]=1;map[216]=0;map[217]=1;map[218]=0;map[219]=1;map[220]=0;
        map[221]=0;map[222]=1;map[223]=1;map[224]=1;map[225]=0;map[226]=1;map[227]=0;map[228]=1;map[229]=0;map[230]=1;map[231]=1;map[232]=1;map[233]=0;map[234]=1;map[235]=0;map[236]=1;map[237]=0;
        map[238]=0;map[239]=1;map[240]=0;map[241]=1;map[242]=0;map[243]=0;map[244]=0;map[245]=0;map[246]=0;map[247]=1;map[248]=0;map[249]=0;map[250]=0;map[251]=0;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=0;map[260]=1;map[261]=1;map[262]=1;map[263]=1;map[264]=1;map[265]=1;map[266]=1;map[267]=0;map[268]=1;map[269]=1;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 5&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=1;map[ 32]=1;map[ 33]=1;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=0;map[ 54]=0;map[ 55]=1;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=0;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=0;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=1;map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=1;map[104]=1;map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=1;map[110]=1;map[111]=0;map[112]=1;map[113]=0;
        map[114]=0;map[115]=1;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;map[121]=1;map[122]=0;map[123]=0;map[124]=0;map[125]=1;map[126]=0;map[127]=1;map[128]=0;map[129]=0;map[130]=0;map[131]=0;map[132]=0;
        map[133]=0;map[134]=1;map[135]=1;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=0;map[142]=1;map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=1;map[148]=1;map[149]=1;map[150]=1;map[151]=0;
        map[152]=0;map[153]=0;map[154]=0;map[155]=1;map[156]=0;map[157]=1;map[158]=0;map[159]=1;map[160]=0;map[161]=1;map[162]=0;map[163]=1;map[164]=0;map[165]=1;map[166]=0;map[167]=0;map[168]=0;map[169]=1;map[170]=0;
        map[171]=0;map[172]=1;map[173]=1;map[174]=1;map[175]=0;map[176]=1;map[177]=0;map[178]=1;map[179]=0;map[180]=1;map[181]=1;map[182]=1;map[183]=0;map[184]=1;map[185]=1;map[186]=1;map[187]=0;map[188]=1;map[189]=0;
        map[190]=0;map[191]=1;map[192]=0;map[193]=1;map[194]=0;map[195]=0;map[196]=0;map[197]=1;map[198]=0;map[199]=0;map[200]=0;map[201]=1;map[202]=0;map[203]=0;map[204]=0;map[205]=0;map[206]=0;map[207]=1;map[208]=0;
        map[209]=0;map[210]=1;map[211]=0;map[212]=1;map[213]=0;map[214]=1;map[215]=1;map[216]=1;map[217]=0;map[218]=1;map[219]=0;map[220]=1;map[221]=1;map[222]=1;map[223]=0;map[224]=1;map[225]=1;map[226]=1;map[227]=0;
        map[228]=0;map[229]=0;map[230]=0;map[231]=0;map[232]=0;map[233]=1;map[234]=0;map[235]=0;map[236]=0;map[237]=1;map[238]=0;map[239]=0;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=0;map[246]=0;
        map[247]=0;map[248]=1;map[249]=1;map[250]=1;map[251]=0;map[252]=1;map[253]=1;map[254]=1;map[255]=0;map[256]=1;map[257]=1;map[258]=1;map[259]=1;map[260]=1;map[261]=0;map[262]=1;map[263]=1;map[264]=1;map[265]=0;
        map[266]=0;map[267]=0;map[268]=0;map[269]=1;map[270]=0;map[271]=1;map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=1;map[278]=0;map[279]=0;map[280]=0;map[281]=1;map[282]=0;map[283]=0;map[284]=0;
        map[285]=0;map[286]=1;map[287]=1;map[288]=1;map[289]=1;map[290]=1;map[291]=0;map[292]=0;map[293]=0;map[294]=1;map[295]=1;map[296]=1;map[297]=1;map[298]=1;map[299]=0;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=0;map[306]=0;map[307]=1;map[308]=0;map[309]=0;map[310]=0;map[311]=1;map[312]=0;map[313]=1;map[314]=0;map[315]=1;map[316]=0;map[317]=1;map[318]=0;map[319]=1;map[320]=0;map[321]=0;map[322]=0;
        map[323]=0;map[324]=1;map[325]=1;map[326]=1;map[327]=0;map[328]=1;map[329]=1;map[330]=1;map[331]=1;map[332]=1;map[333]=0;map[334]=1;map[335]=0;map[336]=1;map[337]=0;map[338]=1;map[339]=1;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 6&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 6&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=1;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=1;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=0;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=0;map[ 32]=0;map[ 33]=0;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=1;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 6&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=1;map[ 60]=0;map[ 61]=0;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=1;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 6&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=1;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=1;map[ 50]=0;map[ 51]=0;map[ 52]=0;map[ 53]=0;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=1;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=1;map[ 74]=0;map[ 75]=1;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=0;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=0;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=0;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=0;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=0;map[104]=1;map[105]=1;map[106]=1;map[107]=1;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;

    end
    if(level == 6&& num == 13)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;
        map[ 13]=0;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=0;
        map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;
        map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;map[ 44]=1;map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=0;map[ 50]=1;map[ 51]=0;
        map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=0;map[ 56]=0;map[ 57]=0;map[ 58]=0;map[ 59]=0;map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=1;map[ 64]=0;
        map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=1;map[ 74]=1;map[ 75]=0;map[ 76]=1;map[ 77]=0;
        map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=0;map[ 88]=0;map[ 89]=1;map[ 90]=0;
        map[ 91]=0;map[ 92]=1;map[ 93]=0;map[ 94]=1;map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=1;map[100]=1;map[101]=0;map[102]=1;map[103]=0;
        map[104]=0;map[105]=0;map[106]=0;map[107]=1;map[108]=0;map[109]=1;map[110]=0;map[111]=1;map[112]=0;map[113]=0;map[114]=0;map[115]=1;map[116]=0;
        map[117]=0;map[118]=1;map[119]=1;map[120]=1;map[121]=0;map[122]=1;map[123]=0;map[124]=1;map[125]=1;map[126]=1;map[127]=0;map[128]=1;map[129]=0;
        map[130]=0;map[131]=1;map[132]=0;map[133]=0;map[134]=0;map[135]=0;map[136]=0;map[137]=1;map[138]=0;map[139]=1;map[140]=0;map[141]=1;map[142]=0;
        map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=1;map[148]=1;map[149]=1;map[150]=1;map[151]=0;map[152]=1;map[153]=0;map[154]=1;map[155]=0;
        map[156]=0;map[157]=0;map[158]=0;map[159]=0;map[160]=0;map[161]=0;map[162]=0;map[163]=0;map[164]=0;map[165]=0;map[166]=0;map[167]=0;map[168]=0;

    end
    if(level == 6&& num == 15)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=0;map[ 20]=1;map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=0;
        map[ 30]=0;map[ 31]=1;map[ 32]=0;map[ 33]=1;map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=1;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=0;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;
        map[ 60]=0;map[ 61]=1;map[ 62]=0;map[ 63]=0;map[ 64]=0;map[ 65]=1;map[ 66]=0;map[ 67]=0;map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=0;map[ 72]=0;map[ 73]=1;map[ 74]=0;
        map[ 75]=0;map[ 76]=1;map[ 77]=0;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=0;map[ 86]=1;map[ 87]=1;map[ 88]=1;map[ 89]=0;
        map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=0;map[ 94]=0;map[ 95]=0;map[ 96]=0;map[ 97]=0;map[ 98]=0;map[ 99]=1;map[100]=0;map[101]=0;map[102]=0;map[103]=1;map[104]=0;
        map[105]=0;map[106]=1;map[107]=1;map[108]=1;map[109]=0;map[110]=1;map[111]=1;map[112]=1;map[113]=1;map[114]=1;map[115]=0;map[116]=1;map[117]=1;map[118]=1;map[119]=0;
        map[120]=0;map[121]=1;map[122]=0;map[123]=0;map[124]=0;map[125]=0;map[126]=0;map[127]=1;map[128]=0;map[129]=1;map[130]=0;map[131]=1;map[132]=0;map[133]=1;map[134]=0;
        map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=1;map[142]=1;map[143]=0;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=0;
        map[150]=0;map[151]=1;map[152]=0;map[153]=0;map[154]=0;map[155]=0;map[156]=0;map[157]=1;map[158]=0;map[159]=1;map[160]=0;map[161]=1;map[162]=0;map[163]=1;map[164]=0;
        map[165]=0;map[166]=1;map[167]=1;map[168]=1;map[169]=0;map[170]=1;map[171]=1;map[172]=1;map[173]=0;map[174]=1;map[175]=0;map[176]=1;map[177]=0;map[178]=1;map[179]=0;
        map[180]=0;map[181]=1;map[182]=0;map[183]=0;map[184]=0;map[185]=0;map[186]=0;map[187]=0;map[188]=0;map[189]=0;map[190]=0;map[191]=0;map[192]=0;map[193]=1;map[194]=0;
        map[195]=0;map[196]=1;map[197]=1;map[198]=1;map[199]=0;map[200]=1;map[201]=1;map[202]=1;map[203]=1;map[204]=1;map[205]=1;map[206]=1;map[207]=1;map[208]=1;map[209]=0;
        map[210]=0;map[211]=0;map[212]=0;map[213]=0;map[214]=0;map[215]=0;map[216]=0;map[217]=0;map[218]=0;map[219]=0;map[220]=0;map[221]=0;map[222]=0;map[223]=0;map[224]=0;

    end
    if(level == 6&& num == 17)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;
        map[ 17]=0;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=0;map[ 32]=0;map[ 33]=0;
        map[ 34]=0;map[ 35]=1;map[ 36]=0;map[ 37]=0;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=1;map[ 50]=0;
        map[ 51]=0;map[ 52]=1;map[ 53]=1;map[ 54]=1;map[ 55]=1;map[ 56]=1;map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=0;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=0;
        map[ 68]=0;map[ 69]=1;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=0;map[ 82]=0;map[ 83]=1;map[ 84]=0;
        map[ 85]=0;map[ 86]=1;map[ 87]=0;map[ 88]=1;map[ 89]=1;map[ 90]=1;map[ 91]=1;map[ 92]=1;map[ 93]=1;map[ 94]=1;map[ 95]=1;map[ 96]=1;map[ 97]=1;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;
        map[102]=0;map[103]=1;map[104]=0;map[105]=1;map[106]=0;map[107]=0;map[108]=0;map[109]=0;map[110]=0;map[111]=0;map[112]=0;map[113]=1;map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;
        map[119]=0;map[120]=1;map[121]=0;map[122]=1;map[123]=1;map[124]=1;map[125]=1;map[126]=1;map[127]=0;map[128]=1;map[129]=1;map[130]=1;map[131]=0;map[132]=1;map[133]=1;map[134]=1;map[135]=0;
        map[136]=0;map[137]=0;map[138]=0;map[139]=1;map[140]=0;map[141]=0;map[142]=0;map[143]=1;map[144]=0;map[145]=0;map[146]=0;map[147]=1;map[148]=0;map[149]=1;map[150]=0;map[151]=0;map[152]=0;
        map[153]=0;map[154]=1;map[155]=1;map[156]=1;map[157]=0;map[158]=1;map[159]=1;map[160]=1;map[161]=0;map[162]=1;map[163]=1;map[164]=1;map[165]=0;map[166]=1;map[167]=1;map[168]=1;map[169]=0;
        map[170]=0;map[171]=0;map[172]=0;map[173]=1;map[174]=0;map[175]=0;map[176]=0;map[177]=0;map[178]=0;map[179]=1;map[180]=0;map[181]=0;map[182]=0;map[183]=1;map[184]=0;map[185]=1;map[186]=0;
        map[187]=0;map[188]=1;map[189]=1;map[190]=1;map[191]=0;map[192]=1;map[193]=1;map[194]=1;map[195]=1;map[196]=1;map[197]=0;map[198]=1;map[199]=1;map[200]=1;map[201]=0;map[202]=1;map[203]=0;
        map[204]=0;map[205]=0;map[206]=0;map[207]=0;map[208]=0;map[209]=1;map[210]=0;map[211]=1;map[212]=0;map[213]=1;map[214]=0;map[215]=0;map[216]=0;map[217]=1;map[218]=0;map[219]=0;map[220]=0;
        map[221]=0;map[222]=1;map[223]=1;map[224]=1;map[225]=1;map[226]=1;map[227]=0;map[228]=1;map[229]=0;map[230]=1;map[231]=0;map[232]=1;map[233]=1;map[234]=1;map[235]=1;map[236]=1;map[237]=0;
        map[238]=0;map[239]=1;map[240]=0;map[241]=1;map[242]=0;map[243]=1;map[244]=0;map[245]=1;map[246]=0;map[247]=0;map[248]=0;map[249]=1;map[250]=0;map[251]=1;map[252]=0;map[253]=1;map[254]=0;
        map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=0;map[260]=1;map[261]=0;map[262]=1;map[263]=0;map[264]=1;map[265]=1;map[266]=1;map[267]=0;map[268]=1;map[269]=0;map[270]=1;map[271]=0;
        map[272]=0;map[273]=0;map[274]=0;map[275]=0;map[276]=0;map[277]=0;map[278]=0;map[279]=0;map[280]=0;map[281]=0;map[282]=0;map[283]=0;map[284]=0;map[285]=0;map[286]=0;map[287]=0;map[288]=0;

    end
    if(level == 6&& num == 19)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;map[ 11]=0;map[ 12]=0;map[ 13]=0;map[ 14]=0;map[ 15]=0;map[ 16]=0;map[ 17]=0;map[ 18]=0;
        map[ 19]=0;map[ 20]=1;map[ 21]=1;map[ 22]=1;map[ 23]=0;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=1;map[ 28]=1;map[ 29]=1;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=1;map[ 36]=1;map[ 37]=0;
        map[ 38]=0;map[ 39]=1;map[ 40]=0;map[ 41]=1;map[ 42]=0;map[ 43]=1;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;map[ 49]=0;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=1;map[ 54]=0;map[ 55]=0;map[ 56]=0;
        map[ 57]=0;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=1;map[ 64]=1;map[ 65]=1;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=1;map[ 72]=1;map[ 73]=0;map[ 74]=1;map[ 75]=0;
        map[ 76]=0;map[ 77]=1;map[ 78]=0;map[ 79]=1;map[ 80]=0;map[ 81]=1;map[ 82]=0;map[ 83]=1;map[ 84]=0;map[ 85]=1;map[ 86]=0;map[ 87]=0;map[ 88]=0;map[ 89]=0;map[ 90]=0;map[ 91]=1;map[ 92]=0;map[ 93]=1;map[ 94]=0;
        map[ 95]=0;map[ 96]=1;map[ 97]=0;map[ 98]=1;map[ 99]=0;map[100]=1;map[101]=0;map[102]=1;map[103]=0;map[104]=1;map[105]=1;map[106]=1;map[107]=1;map[108]=1;map[109]=1;map[110]=1;map[111]=1;map[112]=1;map[113]=0;
        map[114]=0;map[115]=1;map[116]=0;map[117]=1;map[118]=0;map[119]=1;map[120]=0;map[121]=0;map[122]=0;map[123]=1;map[124]=0;map[125]=0;map[126]=0;map[127]=0;map[128]=0;map[129]=0;map[130]=0;map[131]=0;map[132]=0;
        map[133]=0;map[134]=1;map[135]=0;map[136]=1;map[137]=0;map[138]=1;map[139]=1;map[140]=1;map[141]=0;map[142]=1;map[143]=1;map[144]=1;map[145]=0;map[146]=1;map[147]=0;map[148]=1;map[149]=1;map[150]=1;map[151]=0;
        map[152]=0;map[153]=1;map[154]=0;map[155]=1;map[156]=0;map[157]=0;map[158]=0;map[159]=1;map[160]=0;map[161]=1;map[162]=0;map[163]=0;map[164]=0;map[165]=1;map[166]=0;map[167]=1;map[168]=0;map[169]=0;map[170]=0;
        map[171]=0;map[172]=1;map[173]=0;map[174]=1;map[175]=0;map[176]=1;map[177]=1;map[178]=1;map[179]=0;map[180]=1;map[181]=1;map[182]=1;map[183]=1;map[184]=1;map[185]=1;map[186]=1;map[187]=1;map[188]=1;map[189]=0;
        map[190]=0;map[191]=0;map[192]=0;map[193]=1;map[194]=0;map[195]=1;map[196]=0;map[197]=0;map[198]=0;map[199]=1;map[200]=0;map[201]=1;map[202]=0;map[203]=1;map[204]=0;map[205]=0;map[206]=0;map[207]=0;map[208]=0;
        map[209]=0;map[210]=1;map[211]=1;map[212]=1;map[213]=0;map[214]=1;map[215]=0;map[216]=1;map[217]=1;map[218]=1;map[219]=0;map[220]=1;map[221]=0;map[222]=1;map[223]=1;map[224]=1;map[225]=1;map[226]=1;map[227]=0;
        map[228]=0;map[229]=1;map[230]=0;map[231]=1;map[232]=0;map[233]=1;map[234]=0;map[235]=0;map[236]=0;map[237]=1;map[238]=0;map[239]=1;map[240]=0;map[241]=0;map[242]=0;map[243]=1;map[244]=0;map[245]=0;map[246]=0;
        map[247]=0;map[248]=1;map[249]=0;map[250]=1;map[251]=0;map[252]=1;map[253]=0;map[254]=1;map[255]=0;map[256]=1;map[257]=0;map[258]=1;map[259]=0;map[260]=1;map[261]=1;map[262]=1;map[263]=1;map[264]=1;map[265]=0;
        map[266]=0;map[267]=1;map[268]=0;map[269]=0;map[270]=0;map[271]=1;map[272]=0;map[273]=1;map[274]=0;map[275]=0;map[276]=0;map[277]=1;map[278]=0;map[279]=1;map[280]=0;map[281]=1;map[282]=0;map[283]=0;map[284]=0;
        map[285]=0;map[286]=1;map[287]=0;map[288]=1;map[289]=1;map[290]=1;map[291]=1;map[292]=1;map[293]=1;map[294]=1;map[295]=0;map[296]=1;map[297]=0;map[298]=1;map[299]=0;map[300]=1;map[301]=1;map[302]=1;map[303]=0;
        map[304]=0;map[305]=1;map[306]=0;map[307]=0;map[308]=0;map[309]=1;map[310]=0;map[311]=1;map[312]=0;map[313]=1;map[314]=0;map[315]=0;map[316]=0;map[317]=1;map[318]=0;map[319]=1;map[320]=0;map[321]=1;map[322]=0;
        map[323]=0;map[324]=1;map[325]=0;map[326]=1;map[327]=1;map[328]=1;map[329]=0;map[330]=1;map[331]=0;map[332]=1;map[333]=0;map[334]=1;map[335]=1;map[336]=1;map[337]=0;map[338]=1;map[339]=0;map[340]=1;map[341]=0;
        map[342]=0;map[343]=0;map[344]=0;map[345]=0;map[346]=0;map[347]=0;map[348]=0;map[349]=0;map[350]=0;map[351]=0;map[352]=0;map[353]=0;map[354]=0;map[355]=0;map[356]=0;map[357]=0;map[358]=0;map[359]=0;map[360]=0;

    end
    if(level == 7&& num == 5)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;
        map[  5]=0;map[  6]=1;map[  7]=1;map[  8]=1;map[  9]=0;
        map[ 10]=0;map[ 11]=1;map[ 12]=0;map[ 13]=1;map[ 14]=0;
        map[ 15]=0;map[ 16]=1;map[ 17]=0;map[ 18]=1;map[ 19]=0;
        map[ 20]=0;map[ 21]=0;map[ 22]=0;map[ 23]=0;map[ 24]=0;

    end
    if(level == 7&& num == 7)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;
        map[  7]=0;map[  8]=1;map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=0;
        map[ 14]=0;map[ 15]=1;map[ 16]=0;map[ 17]=1;map[ 18]=0;map[ 19]=0;map[ 20]=0;
        map[ 21]=0;map[ 22]=1;map[ 23]=1;map[ 24]=1;map[ 25]=1;map[ 26]=1;map[ 27]=0;
        map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=0;map[ 32]=0;map[ 33]=1;map[ 34]=0;
        map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=1;map[ 40]=1;map[ 41]=0;
        map[ 42]=0;map[ 43]=0;map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=0;map[ 48]=0;

    end
    if(level == 7&& num == 9)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;
        map[  9]=0;map[ 10]=1;map[ 11]=1;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=0;
        map[ 18]=0;map[ 19]=1;map[ 20]=0;map[ 21]=1;map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;
        map[ 27]=0;map[ 28]=1;map[ 29]=0;map[ 30]=1;map[ 31]=0;map[ 32]=1;map[ 33]=0;map[ 34]=1;map[ 35]=0;
        map[ 36]=0;map[ 37]=1;map[ 38]=0;map[ 39]=0;map[ 40]=0;map[ 41]=0;map[ 42]=0;map[ 43]=0;map[ 44]=0;
        map[ 45]=0;map[ 46]=1;map[ 47]=1;map[ 48]=1;map[ 49]=1;map[ 50]=1;map[ 51]=1;map[ 52]=1;map[ 53]=0;
        map[ 54]=0;map[ 55]=1;map[ 56]=0;map[ 57]=1;map[ 58]=0;map[ 59]=0;map[ 60]=0;map[ 61]=1;map[ 62]=0;
        map[ 63]=0;map[ 64]=1;map[ 65]=0;map[ 66]=1;map[ 67]=1;map[ 68]=1;map[ 69]=0;map[ 70]=1;map[ 71]=0;
        map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;map[ 77]=0;map[ 78]=0;map[ 79]=0;map[ 80]=0;

    end
    if(level == 7&& num == 11)begin
        map[  0]=0;map[  1]=0;map[  2]=0;map[  3]=0;map[  4]=0;map[  5]=0;map[  6]=0;map[  7]=0;map[  8]=0;map[  9]=0;map[ 10]=0;
        map[ 11]=0;map[ 12]=1;map[ 13]=1;map[ 14]=1;map[ 15]=1;map[ 16]=1;map[ 17]=1;map[ 18]=1;map[ 19]=1;map[ 20]=1;map[ 21]=0;
        map[ 22]=0;map[ 23]=1;map[ 24]=0;map[ 25]=1;map[ 26]=0;map[ 27]=1;map[ 28]=0;map[ 29]=1;map[ 30]=0;map[ 31]=1;map[ 32]=0;
        map[ 33]=0;map[ 34]=1;map[ 35]=0;map[ 36]=1;map[ 37]=0;map[ 38]=1;map[ 39]=0;map[ 40]=1;map[ 41]=0;map[ 42]=1;map[ 43]=0;
        map[ 44]=0;map[ 45]=0;map[ 46]=0;map[ 47]=1;map[ 48]=0;map[ 49]=0;map[ 50]=0;map[ 51]=1;map[ 52]=0;map[ 53]=1;map[ 54]=0;
        map[ 55]=0;map[ 56]=1;map[ 57]=1;map[ 58]=1;map[ 59]=0;map[ 60]=1;map[ 61]=1;map[ 62]=1;map[ 63]=0;map[ 64]=1;map[ 65]=0;
        map[ 66]=0;map[ 67]=1;map[ 68]=0;map[ 69]=0;map[ 70]=0;map[ 71]=1;map[ 72]=0;map[ 73]=0;map[ 74]=0;map[ 75]=0;map[ 76]=0;
        map[ 77]=0;map[ 78]=1;map[ 79]=1;map[ 80]=1;map[ 81]=0;map[ 82]=1;map[ 83]=1;map[ 84]=1;map[ 85]=1;map[ 86]=1;map[ 87]=0;
        map[ 88]=0;map[ 89]=1;map[ 90]=0;map[ 91]=0;map[ 92]=0;map[ 93]=0;map[ 94]=0;map[ 95]=1;map[ 96]=0;map[ 97]=1;map[ 98]=0;
        map[ 99]=0;map[100]=1;map[101]=1;map[102]=1;map[103]=1;map[104]=1;map[105]=0;map[106]=1;map[107]=0;map[108]=1;map[109]=0;
        map[110]=0;map[111]=0;map[112]=0;map[113]=0;map[114]=0;map[115]=0;map[116]=0;map[117]=0;map[118]=0;map[119]=0;map[120]=0;
    end
    end
end
endmodule